library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

Package MY4 is
	Procedure SQ4(Signal HPOS, VPOS, Points : in integer;
					 Constant MinX, MinY : in integer;
					 Signal DRAW : out std_logic);
End MY4;

Package BODY MY4 is
	Procedure SQ4(Signal HPOS, VPOS, Points : in integer;
					 Constant MinX, MinY : in integer;
					 Signal DRAW : out std_logic) is
					 
	constant letter_s : std_logic_vector(399 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111000000000000010000000000000000000100000000000000000001111111000000000000000000010000000000000000000100000000000000000001000000000000000000010000000000000000000100000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	constant letter_c : std_logic_vector(399 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000110000100000000000011000000000000000000110000000000000000001100000000000000000011000000000000000000110000000000000000001100000000000000000011000001000000000000011111100000000000000000000000000000000000000000000000000000000000000000";
	constant letter_o : std_logic_vector(399 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000011000001100000000001100000001100000000011000000011000000000110000000110000000001100000001100000000011000000011000000000110000000110000000000110000011000000000000011111000000000000000000000000000000000000000000000";
	constant letter_r : std_logic_vector(399 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000000000000011000010000000000000110000110000000000001100001000000000000011111100000000000000110000110000000000001100000110000000000011000000110000000000110000001100000000001100000011000000000000000000000000000000000000000000";
	constant letter_e : std_logic_vector(399 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000110000000000000000001100000000000000000011000000000000000000111110000000000000001111100000000000000011000000000000000000110000000000000000001100000000000000000011111111110000000000000000000000";
	constant letter_ddot : std_logic_vector(399 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000001111000000000000000000000000000";
	
	constant number_0 : std_logic_vector(399 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100000000000011000001100000000001100000001100000000011000000011000000000110000000110000000001100000001100000000011000000011000000000110000000110000000000110000011000000000000111111100000000000000000000000000";
	constant number_1 : std_logic_vector(399 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000011100000000000000001011000000000000000100110000000000000000001100000000000000000011000000000000000000110000000000000000001100000000000000000011000000000000001111111111000000000000000000000000";
	constant number_2 : std_logic_vector(399 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000000000000110000110000000000000000001100000000000000000110000000000000000011000000000000000001100000000000000000110000000000000000011000000000000000011000000000000000001111111111100000000000000000000000";
	constant number_3 : std_logic_vector(399 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000011000000011000000000000000000110000000000000000011000000000000000011100000000000000000001100000000000000000001100000000011000000011000000000001111111000000000000000000000000";
	constant number_4 : std_logic_vector(399 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000001110000000000000000110100000000000000011001000000000000001100010000000000000110000100000000000011000001000000000001111111111100000000000000000100000000000000000001000000000000000000000000";
	constant number_5 : std_logic_vector(399 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000001100000000000000000011000000000000000000011111100000000000000000001100000000000000000001100000000000000000001000000000000000000110000000000001100011000000000000001111100000000000000000000000000";
	
	Begin
			if (HPOS >= (500 + MinX) AND HPOS < (640 + MinX) AND MinY <= VPOS AND VPOS < (20 + MinY)) then
			
				if(HPOS < (520 + MinX)) then
					if(letter_s( ( 399 - ((20 * (VPOS - MinY)) + ((HPOS - MinX) mod 500)) ) ) = '1') then
						DRAW <= '1';
					else
						DRAW <= '0';
					end if;
					
				elsif((520 + MinX) <= HPOS AND HPOS < (540 + MinX)) then
					if(letter_c( ( 399 - ((20 * (VPOS - MinY)) + ((HPOS - MinX) mod 500)) ) ) = '1') then
						DRAW <= '1';
					else
						DRAW <= '0';
					end if; 
					
				elsif((540 + MinX) <= HPOS AND HPOS < (560 + MinX)) then
					if(letter_o( ( 399 - ((20 * (VPOS - MinY)) + ((HPOS - MinX) mod 500)) ) ) = '1') then
						DRAW <= '1';
					else
						DRAW <= '0';
					end if;
					
				elsif((560 + MinX) <= HPOS AND HPOS < (580 + MinX)) then
					if(letter_r( ( 399 - ((20 * (VPOS - MinY)) + ((HPOS - MinX) mod 500)) ) ) = '1') then
						DRAW <= '1';
					else
						DRAW <= '0';
					end if;
					
				elsif((580 + MinX) <= HPOS AND HPOS < (600 + MinX)) then
					if(letter_e( ( 399 - ((20 * (VPOS - MinY)) + ((HPOS - MinX) mod 500)) ) ) = '1') then
						DRAW <= '1';
					else
						DRAW <= '0';
					end if;
					
				elsif((600 + MinX) <= HPOS AND HPOS < (620 + MinX)) then
					if(letter_ddot( ( 399 - ((20 * (VPOS - MinY)) + ((HPOS - MinX) mod 500)) ) ) = '1') then
						DRAW <= '1';
					else
						DRAW <= '0';
					end if;
					
				elsif((620 + MinX) <= HPOS AND HPOS < (640 + MinX)) then
					
					if( Points = 0) then
						if(number_0( ( 399 - ((20 * (VPOS - MinY)) + ((HPOS - MinX) mod 500)) ) ) = '1') then
								DRAW <= '1';
							else
								DRAW <= '0';
							end if;
					end if;
					
					if( Points = 1) then
						if(number_1( ( 399 - ((20 * (VPOS - MinY)) + ((HPOS - MinX) mod 500)) ) ) = '1') then
								DRAW <= '1';
							else
								DRAW <= '0';
							end if;
					end if;
					
					if( Points = 2) then
						if(number_2( ( 399 - ((20 * (VPOS - MinY)) + ((HPOS - MinX) mod 500)) ) ) = '1') then
								DRAW <= '1';
							else
								DRAW <= '0';
							end if;
					end if;
					
					if( Points = 3) then
						if(number_3( ( 399 - ((20 * (VPOS - MinY)) + ((HPOS - MinX) mod 500)) ) ) = '1') then
								DRAW <= '1';
							else
								DRAW <= '0';
							end if;
					end if;
					
					if( Points = 4) then
						if(number_4( ( 399 - ((20 * (VPOS - MinY)) + ((HPOS - MinX) mod 500)) ) ) = '1') then
								DRAW <= '1';
							else
								DRAW <= '0';
							end if;
					end if;
					
					if( Points = 5) then
						if(number_5( ( 399 - ((20 * (VPOS - MinY)) + ((HPOS - MinX) mod 500)) ) ) = '1') then
								DRAW <= '1';
							else
								DRAW <= '0';
							end if;
					end if;
					
					
				end if;
			else
			end if;
			
	end SQ4;
end MY4;